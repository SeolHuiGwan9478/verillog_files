module SYNC_CNT(COUNT,RSTN, CLK, Q0, Q1, Q2);
	input RSTN, CLK, COUNT;
	output Q0, Q1, Q2;

	JK_FF_RESET JK1(Q0,COUNT,COUNT,CLK,RSTN);
	JK_FF_RESET JK2(Q1,Q0,Q0,CLK,RSTN);
	JK_FF_RESET JK3(Q2,(Q1&Q0),(Q1&Q0),CLK,RSTN);

endmodule
		